`define DEPTH 16
`define WIDTH 8
